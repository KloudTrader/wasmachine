`default_nettype none

module fpu64_unary(
  input clk,

  input  [ 2:0] op,
  input  [63:0] a,
  output [63:0] result
);

endmodule
