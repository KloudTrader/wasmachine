`define HAS_MEMORY 0
