`define NONE 0

`define PUSH    1
`define POP     2
`define REPLACE 3

`define EMPTY     1
`define FULL      2
`define UNDERFLOW 3
`define OVERFLOW  4
