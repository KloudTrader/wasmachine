`default_nettype none

module fpu64_binary(
  input clk,

  input  [ 2:0] op,
  input  [63:0] a,
  input  [63:0] b,
  output [63:0] result
);

endmodule
