`default_nettype none

module fpu32;
endmodule
