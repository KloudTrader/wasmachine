`include "stack.vh"

`define UNDERFLOW_RESET       4
`define UNDERFLOW_RESET_PUSH  5
`define UNDERFLOW_GET         6
`define UNDERFLOW_SET         7

`define FULL       4
`define BAD_OFFSET 5
`define BAD_INDEX  6
