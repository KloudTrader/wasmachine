`include "stack.vh"

`define INDEX_RESET 3

`define FULL       4
`define BAD_INDEX  5
