`define i32 2'b00
`define i64 2'b01
`define f32 2'b10
`define f64 2'b11
