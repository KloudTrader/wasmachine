`define NONE 0

`define PUSH    1
`define POP     2
`define REPLACE 3

`define EMPTY     1
`define UNDERFLOW 2
`define OVERFLOW  3
