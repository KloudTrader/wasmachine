`include "stack.vh"

`define INDEX_RESET           4
`define INDEX_RESET_AND_PUSH  5
`define UNDERFLOW_GET         6
`define UNDERFLOW_SET         7

`define FULL       4
`define BAD_OFFSET 5
