`define i32 2'b00
`define i64 2'b01
`define f32 2'b10
`define f64 2'b11

// Traps
`define NONE           0
`define STACK_ERROR    1
`define ROM_ERROR      2
`define UNREACHABLE    3
`define ENDED          4
`define TYPE_MISMATCH  5
`define UNKOWN_OPCODE  6
`define TYPES_MISMATCH 7
