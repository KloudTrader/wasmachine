`include "LimitedStack.vh"

`define REPLACE               4
`define INDEX_RESET_AND_PUSH  5
`define UNDERFLOW_GET         6
`define UNDERFLOW_SET         7

`define BAD_OFFSET 6
